package mem_control_pkg;
    parameter MEM_WIDTH_CODE    = 3;
    parameter mem_lb            = 3'b000;
    parameter mem_lbu           = 3'b001;
    parameter mem_lh            = 3'b010;
    parameter mem_lhu           = 3'b011;
    parameter mem_lw            = 3'b100;
    parameter mem_sb            = 3'b101;
    parameter mem_sh            = 3'b110;
    parameter mem_sw            = 3'b111;
endpackage
